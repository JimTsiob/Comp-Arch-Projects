library verilog;
use verilog.vl_types.all;
entity OR_2_vlg_vec_tst is
end OR_2_vlg_vec_tst;
