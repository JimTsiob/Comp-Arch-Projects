library verilog;
use verilog.vl_types.all;
entity NOT1_vlg_vec_tst is
end NOT1_vlg_vec_tst;
