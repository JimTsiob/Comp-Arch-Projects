LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


ENTITY AND_4 IS 

PORT ( IN1 , IN2, IN3, IN4 : IN STD_LOGIC;
		 OUT1 : OUT STD_LOGIC);
		 
END AND_4;



ARCHITECTURE LOGICFUNC OF AND_4 IS



COMPONENT AND_2 IS 

PORT ( IN1 , IN2 : IN STD_LOGIC;
		 OUT1 : OUT STD_LOGIC);
		 
END COMPONENT;



SIGNAL S1,S2 : STD_LOGIC;

BEGIN 


V0: AND_2 PORT MAP (IN1,IN2,S1);
V1: AND_2 PORT MAP (IN3,IN4,S2);
V2: AND_2 PORT MAP (S1,S2,OUT1);

	
END LOGICFUNC;
