library verilog;
use verilog.vl_types.all;
entity OR_3_vlg_vec_tst is
end OR_3_vlg_vec_tst;
