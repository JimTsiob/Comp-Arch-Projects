library verilog;
use verilog.vl_types.all;
entity NOT1_vlg_sample_tst is
    port(
        A               : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end NOT1_vlg_sample_tst;
