library verilog;
use verilog.vl_types.all;
entity AND_2_vlg_vec_tst is
end AND_2_vlg_vec_tst;
