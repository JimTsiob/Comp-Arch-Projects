library verilog;
use verilog.vl_types.all;
entity XOR_2_vlg_vec_tst is
end XOR_2_vlg_vec_tst;
