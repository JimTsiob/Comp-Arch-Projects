library verilog;
use verilog.vl_types.all;
entity XOR_3 is
    port(
        IN1             : in     vl_logic;
        IN2             : in     vl_logic;
        IN3             : in     vl_logic;
        OUT1            : out    vl_logic
    );
end XOR_3;
