library verilog;
use verilog.vl_types.all;
entity FULLADDER_16_vlg_vec_tst is
end FULLADDER_16_vlg_vec_tst;
