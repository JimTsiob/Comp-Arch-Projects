library verilog;
use verilog.vl_types.all;
entity XOR_3_vlg_check_tst is
    port(
        OUT1            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end XOR_3_vlg_check_tst;
