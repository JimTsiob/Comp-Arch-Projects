library verilog;
use verilog.vl_types.all;
entity OR_3_vlg_check_tst is
    port(
        OUT1            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end OR_3_vlg_check_tst;
