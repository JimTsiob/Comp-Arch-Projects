library verilog;
use verilog.vl_types.all;
entity OR_2 is
    port(
        IN1             : in     vl_logic;
        IN2             : in     vl_logic;
        OUT1            : out    vl_logic
    );
end OR_2;
