library verilog;
use verilog.vl_types.all;
entity XOR_3_vlg_vec_tst is
end XOR_3_vlg_vec_tst;
