library verilog;
use verilog.vl_types.all;
entity AND_2_vlg_check_tst is
    port(
        OUT1            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end AND_2_vlg_check_tst;
