library verilog;
use verilog.vl_types.all;
entity FULLADDER_1_vlg_vec_tst is
end FULLADDER_1_vlg_vec_tst;
