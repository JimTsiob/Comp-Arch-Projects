library verilog;
use verilog.vl_types.all;
entity NOT1 is
    port(
        A               : in     vl_logic;
        Q               : out    vl_logic
    );
end NOT1;
